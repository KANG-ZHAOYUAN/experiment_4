//���������������źţ�ģ��Ľӿڶ������£�

//ģ�����ƣ�key_debounce_15ms
//�����������Ի�е���������źŽ���15ms��ʱ������������ȶ��İ����źż���������/�½�������
//�����źţ�
//  clk      ��ϵͳ�̶�ʱ�ӣ�Ƶ��100MHz
//  rst      ���첽��λ�źţ�����Ч����Ӧʵ����S1������λ������λ�źŲ���Ҫ������������
//  key_in   ��ԭʼ�������루��Ӧʵ����S3����������е������
//����źţ�
//  key_out  ��15ms��ʱ��������ȶ��������
//  rise_pulse�����������������壨1��clk���ڸߵ�ƽ������S3������
//  fall_pulse���������½������壨1��clk���ڸߵ�ƽ�����ã�

module key_debounce_15ms (
    input  wire        clk,         // ϵͳ�̶�ʱ�ӣ�100MHz
    input  wire        rst,         // �첽��λ�źţ�����Ч����Ӧʵ����S1������λ������λ�źŲ���Ҫ������������
    input  wire        key_in,      // ԭʼ�������루��Ӧʵ����S3����������е������
    output reg         key_out,     // 15ms��ʱ��������ȶ��������
    output reg         rise_pulse,  // ���������������壨1��clk���ڸߵ�ƽ������S3������
    output reg         fall_pulse   // �������½������壨1��clk���ڸߵ�ƽ�����ã�
    //rise_pulse��һ�������źţ�ֻ����һ��ʱ��������Ϊ�ߵ�ƽ�����ڴ���S3�����ļ���������
    //fall_pulseҲ��һ�������źţ�ֻ����һ��ʱ��������Ϊ�ߵ�ƽ��ͨ�����ڼ��S3�������ɿ�������
    //��Ȼ�ڱ�ʵ���У�fall_pulse��û��û��ֱ��ʹ�ã�����������Ϊ�����źţ��Ա��������ܵĹ�����չ��
);


parameter DEBOUNCE_CNT_MAX = 21'd1_500_000;
//2^21-1 = 2,097,151���㹻����1,500,000  
// 19λ����������0~750000������15ms������
//���㷽����15ms / 10ns = 1,500,000��ʱ�����ڣ�100MHzʱ������Ϊ10ns��

//�ڲ��źŶ���
reg [2:0]  sync_key;         // ������������ͬ���Ĵ�������������̬��ʵ��ʱ���ȶ���Ҫ��
reg [20:0] debounce_cnt;     // 15ms������������21λ��ƥ��DEBOUNCE_CNT_MAX��
reg        prev_key_out;     // ��һ�����ȶ���������ڱ��ؼ�⣩

// -------------------------- ����1����������ͬ������ --------------------------
// �߼���ʹ�������Ĵ����԰��������źŽ���ͬ����
always @(posedge clk or posedge rst) begin
    if (rst) begin
        sync_key[0] <= 1'b0;
        sync_key[1] <= 1'b0;
        sync_key[2] <= 1'b0;
    end else begin
        sync_key[0] <= key_in;      // ��һ��ͬ�����ɼ�S3ԭʼ�ź�
        sync_key[1] <= sync_key[0]; // �ڶ���ͬ�����ȶ�ͬ�����źţ���������̬
        sync_key[2] <= sync_key[1]; // �������Ĵ��������ã������ڽ�һ���ȶ�����Թ۲�
    end
end
//��ʵ����̫��ȫ�ˣ�ʹ�������Ĵ���ͬ�������źţ��źŻ�������ʱ�����ڵ�������߼�


// -------------------------- ����2��15ms���������� --------------------------
// �߼�����ͬ���󰴼���sync_key[1]���뵱ǰ�ȶ������key_out����һ��ʱ������15ms������
// ������750000��15ms����ֹͣ������ȷ�ϰ���������̬��״̬һ��ʱ���������㡣
always @(posedge clk or posedge rst) begin
    if (rst) begin
        debounce_cnt <= 21'd0;
    end else if (sync_key[2] != key_out) begin  // ��⵽S3״̬�仯����������
        if (debounce_cnt < DEBOUNCE_CNT_MAX) begin
            debounce_cnt <= debounce_cnt + 1'b1; // �������������ۼ�15ms
        end else begin
            debounce_cnt <= debounce_cnt;        // ������15ms��������ֵ�ȴ���̬ȷ��
        end
    end else begin                              // S3״̬�ޱ仯���ȶ��򶶶�������
        debounce_cnt <= 21'd0;                  // ���������㣬���µȴ�״̬�仯
        //ֻҪ�ڶ������ͻ�һֱ����
    end
end

// -------------------------- ����3��15ms��ʱ������ȶ���� --------------------------
// �߼�����������750000��15ms��ʱ��ȷ��S3״̬�ȶ�����ͬ�����źŸ�ֵ��key_out
always @(posedge clk or posedge rst) begin
    if (rst) begin
        key_out <= 1'b0; 
    end else if (debounce_cnt == DEBOUNCE_CNT_MAX) begin
        key_out <= sync_key[2];  // 15ms��ʱ��ȷ����̬�������ȶ����
    end else begin
        key_out <= key_out;      // δ�ﵽ15ms������ԭ�ȶ���������˶���
    end
end

// -------------------------- ����4������������/�½������� --------------------------
// �߼����Աȵ�ǰ�ȶ������key_out������һ���������prev_key_out�������S3�ȶ�����
always @(posedge clk or posedge rst) begin
    if (rst) begin
        prev_key_out <= 1'b0;
        rise_pulse   <= 1'b0;
        fall_pulse   <= 1'b0;
        //�ر�ע��fall_pulse�������Ǳ���0����"�����ź��½�"ʱ��fall_pulse��ʵ��������
    end else begin
        prev_key_out <= key_out;  // �洢��ǰ�ȶ������������һ���ڱ��ضԱ�
        // �����أ�S3���ȶ��͡��ȶ��ߣ���Ӧʵ����S3�����¡�����������������
        rise_pulse <= key_out & ~prev_key_out;
        // �½��أ�S3���ȶ��ߡ��ȶ��ͣ���Ӧʵ����S3���ɿ������������ã�
        fall_pulse <= ~key_out & prev_key_out;
    end
end

endmodule